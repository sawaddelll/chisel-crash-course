module ALU( // @[:@3.2]
  input        clock, // @[:@4.4]
  input        reset, // @[:@5.4]
  input  [7:0] io_a_0, // @[:@6.4]
  input  [7:0] io_b_0, // @[:@6.4]
  input  [2:0] io_ctrl, // @[:@6.4]
  output [7:0] io_result_0, // @[:@6.4]
  output       io_negative, // @[:@6.4]
  output       io_zero, // @[:@6.4]
  output       io_overflow // @[:@6.4]
);
  wire  _T_75; // @[Adder.scala 31:20:@14.4]
  wire  _T_76; // @[Adder.scala 33:27:@19.6]
  wire [8:0] _T_77; // @[Adder.scala 34:27:@21.8]
  wire [7:0] _T_78; // @[Adder.scala 34:27:@22.8]
  wire  _T_79; // @[Adder.scala 35:27:@26.8]
  wire [8:0] _T_80; // @[Adder.scala 36:27:@28.10]
  wire [8:0] _T_81; // @[Adder.scala 36:27:@29.10]
  wire [7:0] _T_82; // @[Adder.scala 36:27:@30.10]
  wire  _T_83; // @[Adder.scala 42:27:@34.10]
  wire [7:0] _T_84; // @[Adder.scala 43:27:@36.12]
  wire  _T_85; // @[Adder.scala 44:27:@40.12]
  wire [7:0] _T_86; // @[Adder.scala 45:27:@42.14]
  wire  _T_87; // @[Adder.scala 46:27:@46.14]
  wire [7:0] _T_88; // @[Adder.scala 47:27:@48.16]
  wire [7:0] _GEN_0; // @[Adder.scala 46:36:@47.14]
  wire [7:0] _GEN_1; // @[Adder.scala 44:35:@41.12]
  wire [7:0] _GEN_2; // @[Adder.scala 42:36:@35.10]
  wire [7:0] _GEN_3; // @[Adder.scala 35:41:@27.8]
  wire [7:0] _GEN_4; // @[Adder.scala 33:36:@20.6]
  wire [7:0] out_0; // @[Adder.scala 31:37:@15.4]
  wire  _T_91; // @[Adder.scala 51:39:@54.4]
  wire  zeroVector_0; // @[Adder.scala 51:24:@55.4]
  wire  _T_94; // @[Adder.scala 56:38:@59.4]
  wire  _T_95; // @[Adder.scala 56:62:@60.4]
  wire  _T_96; // @[Adder.scala 56:51:@61.4]
  wire  _T_97; // @[Adder.scala 56:86:@62.4]
  wire  _T_99; // @[Adder.scala 56:99:@64.4]
  wire  _T_102; // @[Adder.scala 61:36:@68.4]
  assign _T_75 = io_ctrl == 3'h0; // @[Adder.scala 31:20:@14.4]
  assign _T_76 = io_ctrl == 3'h1; // @[Adder.scala 33:27:@19.6]
  assign _T_77 = io_a_0 + io_b_0; // @[Adder.scala 34:27:@21.8]
  assign _T_78 = io_a_0 + io_b_0; // @[Adder.scala 34:27:@22.8]
  assign _T_79 = io_ctrl == 3'h2; // @[Adder.scala 35:27:@26.8]
  assign _T_80 = io_a_0 - io_b_0; // @[Adder.scala 36:27:@28.10]
  assign _T_81 = $unsigned(_T_80); // @[Adder.scala 36:27:@29.10]
  assign _T_82 = _T_81[7:0]; // @[Adder.scala 36:27:@30.10]
  assign _T_83 = io_ctrl == 3'h3; // @[Adder.scala 42:27:@34.10]
  assign _T_84 = io_a_0 & io_b_0; // @[Adder.scala 43:27:@36.12]
  assign _T_85 = io_ctrl == 3'h4; // @[Adder.scala 44:27:@40.12]
  assign _T_86 = io_a_0 | io_b_0; // @[Adder.scala 45:27:@42.14]
  assign _T_87 = io_ctrl == 3'h5; // @[Adder.scala 46:27:@46.14]
  assign _T_88 = io_a_0 ^ io_b_0; // @[Adder.scala 47:27:@48.16]
  assign _GEN_0 = _T_87 ? _T_88 : 8'h0; // @[Adder.scala 46:36:@47.14]
  assign _GEN_1 = _T_85 ? _T_86 : _GEN_0; // @[Adder.scala 44:35:@41.12]
  assign _GEN_2 = _T_83 ? _T_84 : _GEN_1; // @[Adder.scala 42:36:@35.10]
  assign _GEN_3 = _T_79 ? _T_82 : _GEN_2; // @[Adder.scala 35:41:@27.8]
  assign _GEN_4 = _T_76 ? _T_78 : _GEN_3; // @[Adder.scala 33:36:@20.6]
  assign out_0 = _T_75 ? io_a_0 : _GEN_4; // @[Adder.scala 31:37:@15.4]
  assign _T_91 = io_result_0 != 8'h0; // @[Adder.scala 51:39:@54.4]
  assign zeroVector_0 = ~ _T_91; // @[Adder.scala 51:24:@55.4]
  assign _T_94 = io_a_0[7]; // @[Adder.scala 56:38:@59.4]
  assign _T_95 = io_b_0[7]; // @[Adder.scala 56:62:@60.4]
  assign _T_96 = _T_94 == _T_95; // @[Adder.scala 56:51:@61.4]
  assign _T_97 = out_0[7]; // @[Adder.scala 56:86:@62.4]
  assign _T_99 = _T_97 != _T_94; // @[Adder.scala 56:99:@64.4]
  assign _T_102 = zeroVector_0 == 1'h0; // @[Adder.scala 61:36:@68.4]
  assign io_result_0 = _T_75 ? io_a_0 : _GEN_4; // @[Adder.scala 60:15:@67.4]
  assign io_negative = io_result_0[7]; // @[Adder.scala 63:17:@77.4]
  assign io_zero = _T_102 == 1'h0; // @[Adder.scala 61:13:@71.4]
  assign io_overflow = _T_96 & _T_99; // @[Adder.scala 62:17:@74.4]
endmodule
